module led( 
  output [3:0] led 
); 

  assign led = 3; 
endmodule 
