module leds( 
  output [3:0] led 
); 

  assign led = 4'b1111; 
endmodule 
