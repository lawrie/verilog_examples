module pc_vga_8x16_80_FF (
	 input		clk,
	 input  [6:0]	ascii_code,
	 input  [3:0]	row,
	 input  [2:0]  col,
	 output wire	row_of_pixels
	 );

RAMB16_S1 BRAM_PC_VGA_0 (
	.CLK(clk),
	.EN(1'b1),
	.WE(1'b0),
	.ADDR({ascii_code[6:1], ~ascii_code[0], row, ~col}),
	.SSR(1'b0),
	.DI(1'b0),
	.DO(row_of_pixels)
	);
	 
  font[7'h40] = 256'h00007c060c3c66c2c0c0c0c2663c00000000000076cccccccccccc0000cc0000;
  font[7'h41] = 256'h000000007cc6c0c0fec67c0030180c000000000076cccccc7c0c78006c381000;
  font[7'h42] = 256'h0000000076cccccc7c0c780000cc00000000000076cccccc7c0c780018306000;
  font[7'h43] = 256'h0000000076cccccc7c0c7800386c38000000003c060c3c666060663c00000000;
  font[7'h44] = 256'h000000007cc6c0c0fec67c006c381000000000007cc6c0c0fec67c0000c60000;
  font[7'h45] = 256'h000000007cc6c0c0fec67c0018306000000000003c1818181818380000660000;
  font[7'h46] = 256'h000000003c18181818183800663c1800000000003c1818181818380018306000;
  font[7'h47] = 256'h00000000c6c6c6fec6c66c381000c60000000000c6c6c6fec6c66c3800386c38;
  font[7'h48] = 256'h00000000fe6660607c6066fe006030180000000077dcd87e1b3b6e0000000000;
  font[7'h49] = 256'h00000000ceccccccccfecccc6c3e0000000000007cc6c6c6c6c67c006c381000;
  font[7'h4A] = 256'h000000007cc6c6c6c6c67c0000c60000000000007cc6c6c6c6c67c0018306000;
  font[7'h4B] = 256'h0000000076cccccccccccc00cc7830000000000076cccccccccccc0018306000;
  font[7'h4C] = 256'h00780c067ec6c6c6c6c6c60000c60000000000007cc6c6c6c6c6c6c67c00c600;
  font[7'h4D] = 256'h000000007cc6c6c6c6c6c6c6c600c6000000000018187ec3c0c0c0c37e181800;
  font[7'h4E] = 256'h00000000fce660606060f060646c380000000000181818ff18ff183c66c30000;
  font[7'h4F] = 256'h00000000f36666666f66627c6666fc00000070d818181818187e1818181b0e00;

  font[7'h50] = 256'h0000000076cccccc7c0c780060301800000000003c1818181818380030180c00;
  font[7'h51] = 256'h000000007cc6c6c6c6c67c00603018000000000076cccccccccccc0060301800;
  font[7'h52] = 256'h00000000666666666666dc00dc76000000000000c6c6c6cedefef6e6c600dc76;
  font[7'h53] = 256'h0000000000000000007e003e6c6c3c000000000000000000007c00386c6c3800;
  font[7'h54] = 256'h000000007cc6c6c060303000303000000000000000c0c0c0c0fe000000000000;
  font[7'h55] = 256'h000000000006060606fe00000000000000001f0c069bce603018ccc6c2c0c000;
  font[7'h56] = 256'h000006063e96ce663018ccc6c2c0c00000000000183c3c3c1818180018180000;
  font[7'h57] = 256'h000000000000366cd86c360000000000000000000000d86c366cd80000000000;
  font[7'h58] = 256'h44114411441144114411441144114411aa55aa55aa55aa55aa55aa55aa55aa55;
  font[7'h59] = 256'h77dd77dd77dd77dd77dd77dd77dd77dd18181818181818181818181818181818;
  font[7'h5A] = 256'h1818181818181818f8181818181818181818181818181818f818f81818181818;
  font[7'h5B] = 256'h3636363636363636f6363636363636363636363636363636fe00000000000000;
  font[7'h5C] = 256'h1818181818181818f818f800000000003636363636363636f606f63636363636;
  font[7'h5D] = 256'h363636363636363636363636363636363636363636363636f606fe0000000000;
  font[7'h5E] = 256'h0000000000000000fe06f636363636360000000000000000fe36363636363636;
  font[7'h5F] = 256'h0000000000000000f818f818181818181818181818181818f800000000000000;

  font[7'h60] = 256'h00000000000000001f181818181818180000000000000000ff18181818181818;
  font[7'h61] = 256'h1818181818181818ff0000000000000018181818181818181f18181818181818;
  font[7'h62] = 256'h0000000000000000ff000000000000001818181818181818ff18181818181818;
  font[7'h63] = 256'h18181818181818181f181f181818181836363636363636363736363636363636;
  font[7'h64] = 256'h00000000000000003f30373636363636363636363636363637303f0000000000;
  font[7'h65] = 256'h0000000000000000ff00f736363636363636363636363636f700ff0000000000;
  font[7'h66] = 256'h363636363636363637303736363636360000000000000000ff00ff0000000000;
  font[7'h67] = 256'h3636363636363636f700f736363636360000000000000000ff00ff1818181818;
  font[7'h68] = 256'h0000000000000000ff363636363636361818181818181818ff00ff0000000000;
  font[7'h69] = 256'h3636363636363636ff0000000000000000000000000000003f36363636363636;
  font[7'h6A] = 256'h00000000000000001f181f181818181818181818181818181f181f0000000000;
  font[7'h6B] = 256'h36363636363636363f000000000000003636363636363636ff36363636363636;
  font[7'h6C] = 256'h1818181818181818ff18ff18181818180000000000000000f818181818181818;
  font[7'h6D] = 256'h18181818181818181f00000000000000ffffffffffffffffffffffffffffffff;
  font[7'h6E] = 256'hffffffffffffffffff00000000000000f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0;
  font[7'h6F] = 256'h0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f000000000000000000ffffffffffffff;

  font[7'h70] = 256'h0000000076dcd8d8d8dc76000000000000000000ccc6c6c6ccd8cccccc780000;
  font[7'h71] = 256'h00000000c0c0c0c0c0c0c0c6c6fe0000000000006c6c6c6c6c6c6cfe00000000;
  font[7'h72] = 256'h00000000fec66030183060c6fe0000000000000070d8d8d8d8d87e0000000000;
  font[7'h73] = 256'h000000c060607c66666666660000000000000000181818181818dc7600000000;
  font[7'h74] = 256'h000000007e183c6666663c187e00000000000000386cc6c6fec6c66c38000000;
  font[7'h75] = 256'h00000000ee6c6c6c6cc6c6c66c380000000000003c666666663e0c18301e0000;
  font[7'h76] = 256'h0000000000007edbdbdb7e000000000000000000c0607ef3dbdb7e0603000000;
  font[7'h77] = 256'h000000001c306060607c6060301c000000000000c6c6c6c6c6c6c6c67c000000;
  font[7'h78] = 256'h0000000000fe0000fe0000fe0000000000000000ff000018187e181800000000;
  font[7'h79] = 256'h000000007e0030180c060c1830000000000000007e000c18306030180c000000;
  font[7'h7A] = 256'h181818181818181818181b1b1b0e00000000000070d8d8d81818181818181818;
  font[7'h7B] = 256'h00000000001818007e00181800000000000000000000dc7600dc760000000000;
  font[7'h7C] = 256'h0000000000000000000000386c6c380000000000000000181800000000000000;
  font[7'h7D] = 256'h00000000000000180000000000000000000000001c3c6c6cec0c0c0c0c0c0f00;
  font[7'h7E] = 256'h0000000000000000006c6c6c6c6cd800000000000000000000f8c86030d87000;
  font[7'h7F] = 256'h00000000007c7c7c7c7c7c7c0000000000000000000000000000000000000000;
	 
endmodule
