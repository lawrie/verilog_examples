module leds(
  output [7:0] leds
); 

  assign leds = 8'b11111111; 

endmodule
